library verilog;
use verilog.vl_types.all;
entity LineMemory_vlg_vec_tst is
end LineMemory_vlg_vec_tst;
