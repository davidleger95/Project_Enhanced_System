library verilog;
use verilog.vl_types.all;
entity LineMemory_vlg_check_tst is
    port(
        hit             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end LineMemory_vlg_check_tst;
