-- cache.vhd

-- Generated using ACDS version 14.0 209 at 2016.02.12.14:39:05

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cache is
	port (
		clk           : in    std_logic                     := '0';             --                clk.clk
		reset         : in    std_logic                     := '0';             --              reset.reset
		SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => '0'); -- external_interface.DQ
		SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    --                   .ADDR
		SRAM_LB_N     : out   std_logic;                                        --                   .LB_N
		SRAM_UB_N     : out   std_logic;                                        --                   .UB_N
		SRAM_CE_N     : out   std_logic;                                        --                   .CE_N
		SRAM_OE_N     : out   std_logic;                                        --                   .OE_N
		SRAM_WE_N     : out   std_logic;                                        --                   .WE_N
		address       : in    std_logic_vector(19 downto 0) := (others => '0'); --  avalon_sram_slave.address
		byteenable    : in    std_logic_vector(1 downto 0)  := (others => '0'); --                   .byteenable
		read          : in    std_logic                     := '0';             --                   .read
		write         : in    std_logic                     := '0';             --                   .write
		writedata     : in    std_logic_vector(15 downto 0) := (others => '0'); --                   .writedata
		readdata      : out   std_logic_vector(15 downto 0);                    --                   .readdata
		readdatavalid : out   std_logic                                         --                   .readdatavalid
	);
end entity cache;

architecture rtl of cache is
	component cache_sram_0 is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(11 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(11 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component cache_sram_0;

begin
				-- David: Commented this stuff out because it was causing errors
				--signal tag <= address(11 downto 5);
				--signal line_0 <= address(4 downto 2);
				--signal word <= address(1 downto 0);
				
				--type cache_type is array (0 to 8) of std_logic_vector(3 downto 0) of std_logic_vector(15 downto 0);
				--signal temp_cache: cache_type;
	sram_0 : component cache_sram_0
		port map (
			clk           => clk,           --                clk.clk
			reset         => reset,         --              reset.reset
			SRAM_DQ       => SRAM_DQ,       -- external_interface.export
			SRAM_ADDR     => SRAM_ADDR,     --                   .export
			SRAM_LB_N     => SRAM_LB_N,     --                   .export
			SRAM_UB_N     => SRAM_UB_N,     --                   .export
			SRAM_CE_N     => SRAM_CE_N,     --                   .export
			SRAM_OE_N     => SRAM_OE_N,     --                   .export
			SRAM_WE_N     => SRAM_WE_N,     --                   .export
			address       => address,       --  avalon_sram_slave.address
			byteenable    => byteenable,    --                   .byteenable
			read          => read,          --                   .read
			write         => write,         --                   .write
			writedata     => writedata,     --                   .writedata
			readdata      => readdata,      --                   .readdata
			readdatavalid => readdatavalid  --                   .readdatavalid
		);
		readOut: process(clk, reset, address)	-- David: removed 'readdata' from process; was causing error
		begin 
			if rising_edge(clk) then
				-- David: is this to change the clock speed, or something different?
				-- Also, I just completed the if statement for proper syntax
				if (0 = 0) then
					
				end if;
				
			end if;
				
			
		end process; 

end architecture rtl; -- of cache
